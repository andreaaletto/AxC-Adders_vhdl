/home/andrea/vhdl_adders/Src/DCT/DCT2D/BAS09.vhd