/home/andrea/vhdl_adders/Src/DCT/DCT2D/BAS11.vhd