/home/andrea/vhdl_adders/Src/Wrappers/PEA14Wrapper.vhd