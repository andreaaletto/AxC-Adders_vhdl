/home/andrea/vhdl_adders/Src/Wrappers/BAS11Wrapper.vhd