/home/andrea/vhdl_adders/Src/DCT/DCT1D/BC121D.vhd