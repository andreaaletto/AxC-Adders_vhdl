/home/andrea/vhdl_adders/Src/Cells/InAx2.vhd