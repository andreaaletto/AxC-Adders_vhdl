/home/andrea/vhdl_adders/Src/Cells/AMA4.vhd