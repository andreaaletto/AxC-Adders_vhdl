/home/andrea/vhdl_adders/Src/Adders/RippleCarry.vhd