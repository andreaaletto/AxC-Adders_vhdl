/home/andrea/vhdl_adders/Src/Wrappers/BC12Wrapper.vhd