/home/andrea/vhdl_adders/Src/Cells/AMA1.vhd