/home/andrea/vhdl_adders/Src/Wrappers/BAS09Wrapper.vhd