/home/andrea/vhdl_adders/Src/DCT/DCT2D/BC12.vhd