/home/andrea/vhdl_adders/Src/DCT/DCT2D/PEA12.vhd