/home/andrea/vhdl_adders/Src/DCT/DCT2D/BAS08.vhd