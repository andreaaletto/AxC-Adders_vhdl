/home/andrea/vhdl_adders/Src/DCT/DCT1D/BAS081D.vhd