/home/andrea/vhdl_adders/Src/Cells/InAx1.vhd