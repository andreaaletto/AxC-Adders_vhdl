/home/andrea/vhdl_adders/Src/Cells/AXA1.vhd