/home/andrea/vhdl_adders/Src/Cells/AXA2.vhd