/home/andrea/vhdl_adders/Src/Wrappers/CB11Wrapper.vhd