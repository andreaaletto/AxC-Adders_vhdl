/home/andrea/vhdl_adders/Src/Cells/AMA3.vhd