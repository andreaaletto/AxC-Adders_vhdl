/home/andrea/vhdl_adders/Src/Common/Packages.vhd