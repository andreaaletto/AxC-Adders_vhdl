/home/andrea/vhdl_adders/Src/Cells/AMA2.vhd