/home/andrea/vhdl_adders/Src/Common/GenericRegister.vhd