/home/andrea/vhdl_adders/Src/Wrappers/BAS08Wrapper.vhd