/home/andrea/vhdl_adders/Src/Wrappers/PEA12Wrapper.vhd