/home/andrea/vhdl_adders/Src/DCT/DCT1D/PEA121D.vhd