/home/andrea/vhdl_adders/Src/DCT/DCT1D/BAS091D.vhd