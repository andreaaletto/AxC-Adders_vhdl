/home/andrea/vhdl_adders/Src/DCT/DCT2D/CB11.vhd