/home/andrea/vhdl_adders/Src/Cells/AXA3.vhd