/home/andrea/vhdl_adders/Src/Cells/FullAdder.vhd