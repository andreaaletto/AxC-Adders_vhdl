/home/andrea/vhdl_adders/Src/DCT/DCT2D/PEA14.vhd