/home/andrea/vhdl_adders/Src/Adders/generic_adder_subtractor.vhd