/home/andrea/vhdl_adders/Src/Cells/InAx3.vhd