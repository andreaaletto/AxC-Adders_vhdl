/home/andrea/vhdl_adders/Src/DCT/DCT1D/CB111D.vhd