/home/andrea/vhdl_adders/Src/DCT/DCT1D/PEA141D.vhd